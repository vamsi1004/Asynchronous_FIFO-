package fifo_pkg;
`include "uvm_pkg.sv"
`include "uvm_macros.svh"
`include "wr_seq_item.sv"
`include "rd_seq_item.sv"
`include "fifo_wr_sequencer.sv"
`include "fifo_rd_sequencer.sv"
`include "wr_sequence.sv"
`include "rd_sequence.sv"
`include "virtual_sequencer.sv"
`include "virtual_sequence.sv"
`include "fifo_wr_driver.sv"
`include "fifo_rd_driver.sv"
`include "fifo_wr_monitor.sv"
`include "fifo_rd_monitor.sv"
`include "fifo_wr_agent.sv"
`include "fifo_rd_agent.sv"
`include "fifo_scoreboard.sv"
`include "fifo_subscriber.sv"
`include "fifo_environment.sv"
`include "fifo_test.sv"
endpackage
